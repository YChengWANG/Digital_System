// testrom.v
// 
// A purely combinational ROM used to generate test cases for EEC 180
// Lab 3.
//

module testrom (
   input [3:0] addr,
   output reg [127:0] data
   );

   always @(*) begin
      // Test 0: match. 0 c
      // Test 1: match. 4 8
      // Test 2: match. 3 b
      // Test 3: match. 2 d
      // Test 4: match. 0 b
      // Test 5: match. 0 a
      // Test 6: match. 0 b
      // Test 7: match. 2 6
      // Test 8: match. 8 b
      // Test 9: match. 3 6
      // Test 10: match. b f
      // Test 11: match. c d
      // Test 12: match. 6 d
      // Test 13: match. 4 6
      // Test 14: match. 6 7
      // Test 15: no match
      case (addr)
         4'b0000: data[7:0] = 8'b10111001;
         4'b0001: data[7:0] = 8'b00010101;
         4'b0010: data[7:0] = 8'b00110101;
         4'b0011: data[7:0] = 8'b00011010;
         4'b0100: data[7:0] = 8'b01111110;
         4'b0101: data[7:0] = 8'b10111100;
         4'b0110: data[7:0] = 8'b01110011;
         4'b0111: data[7:0] = 8'b01111011;
         4'b1000: data[7:0] = 8'b01001000;
         4'b1001: data[7:0] = 8'b10100010;
         4'b1010: data[7:0] = 8'b11100001;
         4'b1011: data[7:0] = 8'b11000010;
         4'b1100: data[7:0] = 8'b10111101;
         4'b1101: data[7:0] = 8'b11111110;
         4'b1110: data[7:0] = 8'b01111111;
         default: data[7:0] = 8'b01000001;
      endcase
      case (addr)
         4'b0000: data[15:8] = 8'b01101000;
         4'b0001: data[15:8] = 8'b11001001;
         4'b0010: data[15:8] = 8'b00101101;
         4'b0011: data[15:8] = 8'b00001101;
         4'b0100: data[15:8] = 8'b00001110;
         4'b0101: data[15:8] = 8'b00011000;
         4'b0110: data[15:8] = 8'b10111010;
         4'b0111: data[15:8] = 8'b01110011;
         4'b1000: data[15:8] = 8'b11011101;
         4'b1001: data[15:8] = 8'b01100011;
         4'b1010: data[15:8] = 8'b00100111;
         4'b1011: data[15:8] = 8'b11101001;
         4'b1100: data[15:8] = 8'b11110110;
         4'b1101: data[15:8] = 8'b11001001;
         4'b1110: data[15:8] = 8'b00000101;
         default: data[15:8] = 8'b10101000;
      endcase
      case (addr)
         4'b0000: data[23:16] = 8'b10110111;
         4'b0001: data[23:16] = 8'b01101100;
         4'b0010: data[23:16] = 8'b10101000;
         4'b0011: data[23:16] = 8'b01000010;
         4'b0100: data[23:16] = 8'b10010001;
         4'b0101: data[23:16] = 8'b11000010;
         4'b0110: data[23:16] = 8'b11100011;
         4'b0111: data[23:16] = 8'b01110000;
         4'b1000: data[23:16] = 8'b00000000;
         4'b1001: data[23:16] = 8'b01100010;
         4'b1010: data[23:16] = 8'b11110001;
         4'b1011: data[23:16] = 8'b10010111;
         4'b1100: data[23:16] = 8'b00101101;
         4'b1101: data[23:16] = 8'b10110101;
         4'b1110: data[23:16] = 8'b01111110;
         default: data[23:16] = 8'b01010111;
      endcase
      case (addr)
         4'b0000: data[31:24] = 8'b11010001;
         4'b0001: data[31:24] = 8'b00110110;
         4'b0010: data[31:24] = 8'b01001000;
         4'b0011: data[31:24] = 8'b00001000;
         4'b0100: data[31:24] = 8'b01001010;
         4'b0101: data[31:24] = 8'b01000100;
         4'b0110: data[31:24] = 8'b00001000;
         4'b0111: data[31:24] = 8'b11100001;
         4'b1000: data[31:24] = 8'b00101011;
         4'b1001: data[31:24] = 8'b10011100;
         4'b1010: data[31:24] = 8'b00100110;
         4'b1011: data[31:24] = 8'b00011101;
         4'b1100: data[31:24] = 8'b10101011;
         4'b1101: data[31:24] = 8'b10101010;
         4'b1110: data[31:24] = 8'b01001111;
         default: data[31:24] = 8'b01100011;
      endcase
      case (addr)
         4'b0000: data[39:32] = 8'b01011011;
         4'b0001: data[39:32] = 8'b01100001;
         4'b0010: data[39:32] = 8'b10011011;
         4'b0011: data[39:32] = 8'b11001001;
         4'b0100: data[39:32] = 8'b01110111;
         4'b0101: data[39:32] = 8'b11111110;
         4'b0110: data[39:32] = 8'b10101100;
         4'b0111: data[39:32] = 8'b11011011;
         4'b1000: data[39:32] = 8'b00010100;
         4'b1001: data[39:32] = 8'b01111110;
         4'b1010: data[39:32] = 8'b11111110;
         4'b1011: data[39:32] = 8'b01000110;
         4'b1100: data[39:32] = 8'b11101001;
         4'b1101: data[39:32] = 8'b00101010;
         4'b1110: data[39:32] = 8'b10110100;
         default: data[39:32] = 8'b01101001;
      endcase
      case (addr)
         4'b0000: data[47:40] = 8'b01110000;
         4'b0001: data[47:40] = 8'b10010001;
         4'b0010: data[47:40] = 8'b01111101;
         4'b0011: data[47:40] = 8'b00010000;
         4'b0100: data[47:40] = 8'b11110011;
         4'b0101: data[47:40] = 8'b01110111;
         4'b0110: data[47:40] = 8'b10110110;
         4'b0111: data[47:40] = 8'b11100000;
         4'b1000: data[47:40] = 8'b01101011;
         4'b1001: data[47:40] = 8'b01110111;
         4'b1010: data[47:40] = 8'b01101010;
         4'b1011: data[47:40] = 8'b11101100;
         4'b1100: data[47:40] = 8'b10001110;
         4'b1101: data[47:40] = 8'b00101100;
         4'b1110: data[47:40] = 8'b11011111;
         default: data[47:40] = 8'b10010110;
      endcase
      case (addr)
         4'b0000: data[55:48] = 8'b00111000;
         4'b0001: data[55:48] = 8'b10100010;
         4'b0010: data[55:48] = 8'b01101111;
         4'b0011: data[55:48] = 8'b10111101;
         4'b0100: data[55:48] = 8'b01101110;
         4'b0101: data[55:48] = 8'b00010010;
         4'b0110: data[55:48] = 8'b01011100;
         4'b0111: data[55:48] = 8'b01001011;
         4'b1000: data[55:48] = 8'b10110100;
         4'b1001: data[55:48] = 8'b10011100;
         4'b1010: data[55:48] = 8'b10101011;
         4'b1011: data[55:48] = 8'b01100110;
         4'b1100: data[55:48] = 8'b11111000;
         4'b1101: data[55:48] = 8'b00101101;
         4'b1110: data[55:48] = 8'b11110010;
         default: data[55:48] = 8'b10011100;
      endcase
      case (addr)
         4'b0000: data[63:56] = 8'b01010010;
         4'b0001: data[63:56] = 8'b11110001;
         4'b0010: data[63:56] = 8'b00101010;
         4'b0011: data[63:56] = 8'b11110001;
         4'b0100: data[63:56] = 8'b01100110;
         4'b0101: data[63:56] = 8'b11110100;
         4'b0110: data[63:56] = 8'b11110010;
         4'b0111: data[63:56] = 8'b10101110;
         4'b1000: data[63:56] = 8'b01011100;
         4'b1001: data[63:56] = 8'b01001111;
         4'b1010: data[63:56] = 8'b11111000;
         4'b1011: data[63:56] = 8'b00000101;
         4'b1100: data[63:56] = 8'b00110100;
         4'b1101: data[63:56] = 8'b01001110;
         4'b1110: data[63:56] = 8'b11110010;
         default: data[63:56] = 8'b01101101;
      endcase
      case (addr)
         4'b0000: data[71:64] = 8'b00010111;
         4'b0001: data[71:64] = 8'b01011111;
         4'b0010: data[71:64] = 8'b11101111;
         4'b0011: data[71:64] = 8'b11101000;
         4'b0100: data[71:64] = 8'b01011010;
         4'b0101: data[71:64] = 8'b01110001;
         4'b0110: data[71:64] = 8'b00010101;
         4'b0111: data[71:64] = 8'b01110000;
         4'b1000: data[71:64] = 8'b01101110;
         4'b1001: data[71:64] = 8'b01000011;
         4'b1010: data[71:64] = 8'b10000101;
         4'b1011: data[71:64] = 8'b11011011;
         4'b1100: data[71:64] = 8'b00111110;
         4'b1101: data[71:64] = 8'b01100111;
         4'b1110: data[71:64] = 8'b11011101;
         default: data[71:64] = 8'b10000101;
      endcase
      case (addr)
         4'b0000: data[79:72] = 8'b11110011;
         4'b0001: data[79:72] = 8'b00100011;
         4'b0010: data[79:72] = 8'b10001111;
         4'b0011: data[79:72] = 8'b01001111;
         4'b0100: data[79:72] = 8'b10000101;
         4'b0101: data[79:72] = 8'b00001001;
         4'b0110: data[79:72] = 8'b11000101;
         4'b0111: data[79:72] = 8'b11111100;
         4'b1000: data[79:72] = 8'b00011011;
         4'b1001: data[79:72] = 8'b00011010;
         4'b1010: data[79:72] = 8'b00001001;
         4'b1011: data[79:72] = 8'b00010001;
         4'b1100: data[79:72] = 8'b10101110;
         4'b1101: data[79:72] = 8'b10101011;
         4'b1110: data[79:72] = 8'b11111100;
         default: data[79:72] = 8'b10111010;
      endcase
      case (addr)
         4'b0000: data[87:80] = 8'b11111100;
         4'b0001: data[87:80] = 8'b01111110;
         4'b0010: data[87:80] = 8'b00111000;
         4'b0011: data[87:80] = 8'b10010101;
         4'b0100: data[87:80] = 8'b10110101;
         4'b0101: data[87:80] = 8'b10111100;
         4'b0110: data[87:80] = 8'b00100110;
         4'b0111: data[87:80] = 8'b11000100;
         4'b1000: data[87:80] = 8'b00111100;
         4'b1001: data[87:80] = 8'b10001110;
         4'b1010: data[87:80] = 8'b10100110;
         4'b1011: data[87:80] = 8'b00010110;
         4'b1100: data[87:80] = 8'b00111111;
         4'b1101: data[87:80] = 8'b00010110;
         4'b1110: data[87:80] = 8'b00000111;
         default: data[87:80] = 8'b01111010;
      endcase
      case (addr)
         4'b0000: data[95:88] = 8'b00101110;
         4'b0001: data[95:88] = 8'b11100101;
         4'b0010: data[95:88] = 8'b01001000;
         4'b0011: data[95:88] = 8'b11010100;
         4'b0100: data[95:88] = 8'b01111110;
         4'b0101: data[95:88] = 8'b00101010;
         4'b0110: data[95:88] = 8'b01110011;
         4'b0111: data[95:88] = 8'b11101000;
         4'b1000: data[95:88] = 8'b01101110;
         4'b1001: data[95:88] = 8'b01000101;
         4'b1010: data[95:88] = 8'b01100101;
         4'b1011: data[95:88] = 8'b00010101;
         4'b1100: data[95:88] = 8'b10101001;
         4'b1101: data[95:88] = 8'b01010010;
         4'b1110: data[95:88] = 8'b10100110;
         default: data[95:88] = 8'b10011010;
      endcase
      case (addr)
         4'b0000: data[103:96] = 8'b10111001;
         4'b0001: data[103:96] = 8'b01100001;
         4'b0010: data[103:96] = 8'b01000001;
         4'b0011: data[103:96] = 8'b00111111;
         4'b0100: data[103:96] = 8'b01001101;
         4'b0101: data[103:96] = 8'b11011001;
         4'b0110: data[103:96] = 8'b11000000;
         4'b0111: data[103:96] = 8'b01001011;
         4'b1000: data[103:96] = 8'b00110100;
         4'b1001: data[103:96] = 8'b11001110;
         4'b1010: data[103:96] = 8'b01011111;
         4'b1011: data[103:96] = 8'b11101011;
         4'b1100: data[103:96] = 8'b10100101;
         4'b1101: data[103:96] = 8'b01001100;
         4'b1110: data[103:96] = 8'b00111101;
         default: data[103:96] = 8'b10100011;
      endcase
      case (addr)
         4'b0000: data[111:104] = 8'b00101010;
         4'b0001: data[111:104] = 8'b01101010;
         4'b0010: data[111:104] = 8'b11100110;
         4'b0011: data[111:104] = 8'b01000010;
         4'b0100: data[111:104] = 8'b11110000;
         4'b0101: data[111:104] = 8'b01011001;
         4'b0110: data[111:104] = 8'b10101001;
         4'b0111: data[111:104] = 8'b10101011;
         4'b1000: data[111:104] = 8'b01110110;
         4'b1001: data[111:104] = 8'b00000000;
         4'b1010: data[111:104] = 8'b01010011;
         4'b1011: data[111:104] = 8'b11101011;
         4'b1100: data[111:104] = 8'b11111000;
         4'b1101: data[111:104] = 8'b00101010;
         4'b1110: data[111:104] = 8'b10100101;
         default: data[111:104] = 8'b11011001;
      endcase
      case (addr)
         4'b0000: data[119:112] = 8'b11010010;
         4'b0001: data[119:112] = 8'b01100110;
         4'b0010: data[119:112] = 8'b01101101;
         4'b0011: data[119:112] = 8'b00000011;
         4'b0100: data[119:112] = 8'b01000110;
         4'b0101: data[119:112] = 8'b11110111;
         4'b0110: data[119:112] = 8'b11011101;
         4'b0111: data[119:112] = 8'b00001111;
         4'b1000: data[119:112] = 8'b00011100;
         4'b1001: data[119:112] = 8'b00101101;
         4'b1010: data[119:112] = 8'b11101110;
         4'b1011: data[119:112] = 8'b01000100;
         4'b1100: data[119:112] = 8'b01001111;
         4'b1101: data[119:112] = 8'b00101101;
         4'b1110: data[119:112] = 8'b01000010;
         default: data[119:112] = 8'b01011011;
      endcase
      case (addr)
         4'b0000: data[127:120] = 8'b10001000;
         4'b0001: data[127:120] = 8'b01011111;
         4'b0010: data[127:120] = 8'b00001000;
         4'b0011: data[127:120] = 8'b10001111;
         4'b0100: data[127:120] = 8'b10101111;
         4'b0101: data[127:120] = 8'b10101011;
         4'b0110: data[127:120] = 8'b11011101;
         4'b0111: data[127:120] = 8'b01011100;
         4'b1000: data[127:120] = 8'b01011010;
         4'b1001: data[127:120] = 8'b01000011;
         4'b1010: data[127:120] = 8'b01100101;
         4'b1011: data[127:120] = 8'b10101011;
         4'b1100: data[127:120] = 8'b11101010;
         4'b1101: data[127:120] = 8'b11010000;
         4'b1110: data[127:120] = 8'b11010110;
         default: data[127:120] = 8'b01110110;
      endcase
   end
endmodule      //testrom