module tb1_compare15;
  wire match; // 0=no match, 1=match
  wire [3:0] num_match_low;
  //output [14:0] kkk;
  reg [7:0] in0, in1, in2, in3, in4, in5, in6, in7,
              in8, in9, ina, inb, inc, ind, ine;
  reg [7:0] cpii;
  reg Enable;
  always@(*)begin
      in0=8'b0000_0000;
	   in1=8'b0000_0000;
	   in2=8'b0000_0000;
	   in3=8'b0000_0000;
	   in4=8'b0000_0000;
	   in5=8'b0000_0000;
	   in6=8'b0000_0000;
	   in7=8'b0000_0000;
	   in8=8'b0000_0000;
	   in9=8'b0000_0000;
	   ina=8'b0000_0000;
	   inb=8'b0000_0000;
	   inc=8'b0000_0000;
	   ind=8'b0000_0000;
	   ine=8'b0000_0000;
	 if(Enable==1)begin
      in0=8'b0000_0001;
	   in1=8'b0000_0010;
	   in2=8'b0000_0100;
	   in3=8'b0000_1000;
	   in4=8'b0001_0000;
	   in5=8'b0010_0000;
	   in6=8'b0100_0000;
	   in7=8'b1000_0000;
	   in8=8'b1000_0001;
	   in9=8'b0100_0010;
	   ina=8'b0010_0100;
	   inb=8'b0001_1000;
	   inc=8'b0110_0110;
	   ind=8'b1001_1001;
	   ine=8'b1111_1111;
	 end
  end	

  compare15 cp1(.compare_input(cpii), .in0(in0), .in1(in1), .in2(in2), 
               .in3(in3), .in4(in4), .in5(in5), .in6(in6), 
               .in7(in7), .in8(in8), .in9(in9), .ina(ina),
               .inb(inb), .inc(inc), .ind(ind), .ine(ine),  
					.match(match), .num_match_low(num_match_low));
				

    initial begin
	  //always@(*)begin
	   Enable=1;
		#100
		cpii=8'b0000_0001;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_0010;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_0100;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_1000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0001_0000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0010_0000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0100_0000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b1000_0000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_0001;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_0010;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_0100;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0000_1000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b1000_0001;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0100_0010;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0010_0100;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0001_1000;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b0110_0110;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b1001_1001;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		#100
		Enable=1;
		#100
		cpii=8'b1111_1111;
		#100
	   $display("%b,%h",match,num_match_low);
      Enable=0;
		$stop;
    //end
	end 
  endmodule